module data_forwarding();

endmodule
